*Full wave Bridge Rectifier
*For 12V RMS, the peak value is 12*1.414 = 16.97V
Vin TxTop TxBottom DC 0 Sin(0 16.97 50 0 0)
D1 TxTop    Out		DF
D2 TxBottom Out		DF
D3 Gnd      TxTop	DF
D4 Gnd	    TxBottom	DF
.MODEL DF D (IS=6.22n N=1.9224 RS=0.336 CJ0=764f VJ=0.75 BV=200 TT=2.88n)

RL Out TestPt 1k
Vtest TestPt Gnd 0V

.tran 100u 60m 20m

.control
run
plot V(TxTop) V(TxBottom)
plot V(TxTop)-V(TxBottom) V(Out)
plot I(Vtest)
.endc
.end

