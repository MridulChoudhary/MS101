*Full wave Bridge Rectifier
*For 12V RMS, the peak value is 12*1.414 = 16.97V
Vin TxTop TxBottom DC 0 Sin(0 16.97 50 0 0)
D1 TxTop    Out		DF
D2 TxBottom Out		DF
D3 Gnd      TxTop	DF
D4 Gnd	    TxBottom	DF
.MODEL DF D (IS=6.22n N=1.9224 RS=0.336 CJ0=764f VJ=0.75 BV=200 TT=2.88n)

RL Out TestPt 500
Vtest TestPt Gnd 0V
C  Out Gnd 100u

.tran 10u 60m

.control
run
plot V(TxTop)- V(TxBottom) V(Out)
plot V(out) ylimit 13.4, 15.8
plot -I(Vin)
.endc
.end

